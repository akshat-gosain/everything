`include "full_adder.v"
module bit4_adder(input [3:0]A,input  [3:0]B,input C0,output  [3:0]O, output C1);
    

endmodule